../chisel/verilog/hb_universal.sv